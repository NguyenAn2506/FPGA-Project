library ieee;
use ieee.std_logic_1164.all;
entity FPGA_LCD_DEM_PC_UART is
	Port(	CKHT	: in 	STD_LOGIC;
			BTN_N0	: in 	STD_LOGIC;
			SW0 	: in 	STD_LOGIC;
			BELL	: out	STD_LOGIC;
			UART_RX	: in 	STD_LOGIC;
			UART_TX	: OUT	STD_LOGIC;
			LCD_E	: OUT	STD_LOGIC;
			LCD_RS	: OUT 	STD_LOGIC;
			LCD_RW	: OUT	STD_LOGIC;
			LCD_DB	: OUT 	STD_LOGIC_VECTOR(7 downto 0)
			);
	END FPGA_LCD_DEM_PC_UART;
	
architecture Behavioral of FPGA_LCD_DEM_PC_UART is
	SIGNAL	RST				: STD_LOGIC;
	SIGNAL	LCD_HANG_1_R	: STD_LOGIC_VECTOR(127 downto 0);
	SIGNAL	LCD_HANG_1_N	: STD_LOGIC_VECTOR(127 downto 0);
	SIGNAL	LCD_HANG_2		: STD_LOGIC_VECTOR(127 downto 0);
			
	SIGNAL	UART_TX_FULL	: STD_LOGIC;
	SIGNAL	UART_RX_EMPTY	: STD_LOGIC;
	
	SIGNAL	UART_RECV_DATA	: STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL	UART_TRANS_DATA	: STD_LOGIC_VECTOR(7 downto 0);
	
	SIGNAL	UART_ENA_TX		: STD_LOGIC;
	SIGNAL 	UART_ENA_RD		: STD_LOGIC;
	
	SIGNAL 	ENA_DB			: STD_LOGIC;
	SIGNAL 	ENA_RX			: STD_LOGIC;
	SIGNAL 	DEM				: STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL 	DONVI 			: STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL 	CHUC 			: STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL 	TRAM 			: STD_LOGIC_VECTOR(3 downto 0);
	
begin
	RST		<= not BTN_N0;
	BELL	<= '1';
	LCD_RW	<= '0';
	ENA_RX	<= CKHT;
	
	CHIA_10ENA	:	ENTITY WORK.CHIA_10ENA
		PORT MAP(	CKHT	=> CKHT,
					ENA5Hz	=> ENA_DB );
	UART_UNIT:	ENTITY WORK.UART_CONTROLLER
		PORT MAP(	CKHT	=> CKHT,
					RST		=> RST,
					UART_RX	=> UART_RX,
					UART_TX	=> UART_TX
					FIFO_UART_RX_ENA_RD		=> UART_ENA_RD,
					FIFO_UART_RX_DATA_RD	=> UART_RECV_DATA,
					FIFO_UART_RX_EMPTY		=> UART_RX_EMPTY,
					FIFO_UART_TX_ENA_WR		=> UART_ENA_TX,
					FIFO_UART_TX_DATA_WR	=> UART_TRANS_DATA,
					FIFO_UART_TX_FULL		=> UART_TX_FULL);
		PROCESS(UART_TX_FULL, ENA_DB, SW0, DEM)
		BEGIN
			UART_TRANS_DATA		<= DEM; 	-- GAN DL DOI DI
			IF	UART_TX_FULL = '0'  THEN
				UART_ENA_TX		<= ENA_DB AND SW0;	-- TAO XUNG PHAT
			ELSE 	
				UART_ENA_TX	<= '0';
			END IF;
		END PROCESS;
		
		UART_ENA_RD		<= ENA_RX AND (NOT UART_RX_EMPTY); 	-- TAO XUNG DOC
		PROCESS(CKHT, RST)
		BEGIN
			IF RST = '1' THEN
				LCD_HANG_1_R <= X"20202020202020202020202020202020";
				ELSIF FALLING_EDGE(CKHT) THEN
					LCD_HANG_1_R <= LCD_HANG_1_N;
			END IF;
		END PROCESS;
		LCD_HANG_1_N <= UART_RECV_DATA & LCD_HANG_1_R(127 downto 8)	
						WHEN UART_ENA_RD = '1'
						ELSE LCD_HANG_1_R;
	
	DEM_8BIT:	ENTITY WORK.DEM_8BIT
		PORT MAP(	CKHT	=> CKHT,
					RST 	=> RST,
					ENA_SS	=> SW0,
					ENA_DB	=> ENA_DB,
					DEM 	=> DEM);
	HEXTOBCD: 	ENTITY WORK.HEXTOBCD_8BIT
		PORT MAP(	SOHEX8BIT	=> DEM,
					DONVI		=> DONVI,
					CHUC		=> CHUC,
					TRAM		=> TRAM);
	LCD_GAN_DULIEU_HIENTHI_H2	: ENTITY WORK.LCD_GAN_DULIEU_HIENTHI_H2
		PORT MAP(	H2_13	=> TRAM,
					H2_14	=> CHUC,
					H2_15	=> DONVI,
					LCD_HANG_2	=> LCD_HANG_2);
	LCD_KHOITAO_HIENTHI: 	ENTITY WORK.LCD_KHOITAO_HIENTHI
		PORT MAP(	LCD_DB	=> LCD_DB,
					LCD_RS	=> LCD_RS,
					LCD_E	=> LCD_E,
					LCD_RST	=> RST,
					LCD_CK	=> CKHT,
					LCD_HANG_1 => LCD_HANG_1_R,
					LCD_HANG_2 => LCD_HANG_2);
END Behavioral;
		
		
		
				
			